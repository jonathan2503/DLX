package CONSTANTS is

   constant ALL_BITS      : integer := 32;	
   constant N_BIT         : integer := 4;	
   constant N_subdiv      : integer := 4;	
   constant N_Block       : integer := 8;	
   constant address_ram   : integer := 16;	
end CONSTANTS;
